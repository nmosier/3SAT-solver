// test if you can read file into parameter

module test();
	localparam file_no fopen("tst/test1.txt");
	
endmodule